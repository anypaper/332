// Copyright (C) 2016
// All rights reserved.
//
//
// @NETFPGA_LICENSE_HEADER_START@
//
// Licensed to NetFPGA C.I.C. (NetFPGA) under one or more contributor
// license agreements.  See the NOTICE file distributed with this work for
// additional information regarding copyright ownership.  NetFPGA licenses this
// file to you under the NetFPGA Hardware-Software License, Version 1.0 (the
// "License"); you may not use this file except in compliance with the
// License.  You may obtain a copy of the License at:
//
//   http://www.netfpga-cic.org
//
// Unless required by applicable law or agreed to in writing, Work distributed
// under the License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied.  See the License for the
// specific language governing permissions and limitations under the License.
//
// @NETFPGA_LICENSE_HEADER_END@
//
/*******************************************************************************
 *  File:
 *        rate_limiter.v
 *
 *  Library:
 *        hw/std/cores/rate_limiter_v1_0_0
 *
 *  Module:
 *        rate_limiter
 *
 *  Author:
 * 		
 *  Description:
 *        rate_limiter module
 *
 */

`timescale 1ns/1ps
`include "rate_limiter_cpu_regs_defines.v"

module rate_limiter
#(
    //Master AXI Stream Data Width
    parameter C_M_AXIS_DATA_WIDTH=512,
    parameter C_S_AXIS_DATA_WIDTH=512,
    parameter C_M_AXIS_TUSER_WIDTH=128,
    parameter C_S_AXIS_TUSER_WIDTH=128,

 // AXI Registers Data Width
    parameter C_S_AXI_DATA_WIDTH    = 32,          
    parameter C_S_AXI_ADDR_WIDTH    = 12,          
    parameter C_BASEADDR            = 32'h00000000


)
(
    // Global Ports
    input axis_aclk,
    input axis_resetn,

    // Master Stream Ports (interface to data path)
    output [C_M_AXIS_DATA_WIDTH - 1:0] m_axis_tdata,
    output [((C_M_AXIS_DATA_WIDTH / 8)) - 1:0] m_axis_tkeep,
    output [C_M_AXIS_TUSER_WIDTH-1:0] m_axis_tuser,
    output m_axis_tvalid,
    input  m_axis_tready,
    output m_axis_tlast,

    // Slave Stream Ports (interface to RX queues)
    input [C_S_AXIS_DATA_WIDTH - 1:0] s_axis_tdata,
    input [((C_S_AXIS_DATA_WIDTH / 8)) - 1:0] s_axis_tkeep,
    input [C_S_AXIS_TUSER_WIDTH-1:0] s_axis_tuser,
    input  s_axis_tvalid,
    output s_axis_tready,
    input  s_axis_tlast,

// Slave AXI Ports
    input                                     S_AXI_ACLK,
    input                                     S_AXI_ARESETN,
    input      [C_S_AXI_ADDR_WIDTH-1 : 0]     S_AXI_AWADDR,
    input                                     S_AXI_AWVALID,
    input      [C_S_AXI_DATA_WIDTH-1 : 0]     S_AXI_WDATA,
    input      [C_S_AXI_DATA_WIDTH/8-1 : 0]   S_AXI_WSTRB,
    input                                     S_AXI_WVALID,
    input                                     S_AXI_BREADY,
    input      [C_S_AXI_ADDR_WIDTH-1 : 0]     S_AXI_ARADDR,
    input                                     S_AXI_ARVALID,
    input                                     S_AXI_RREADY,
    output                                    S_AXI_ARREADY,
    output     [C_S_AXI_DATA_WIDTH-1 : 0]     S_AXI_RDATA,
    output     [1 : 0]                        S_AXI_RRESP,
    output                                    S_AXI_RVALID,
    output                                    S_AXI_WREADY,
    output     [1 :0]                         S_AXI_BRESP,
    output                                    S_AXI_BVALID,
    output                                    S_AXI_AWREADY
);

   reg      [`REG_ID_BITS]    id_reg;
   reg      [`REG_VERSION_BITS]    version_reg;
   wire     [`REG_RESET_BITS]    reset_reg;
   reg      [`REG_FLIP_BITS]    ip2cpu_flip_reg;
   wire     [`REG_FLIP_BITS]    cpu2ip_flip_reg;
   reg      [`REG_PKTIN_BITS]    pktin_reg;
   wire                             pktin_reg_clear;
   reg      [`REG_PKTOUT_BITS]    pktout_reg;
   wire                             pktout_reg_clear;
   reg      [`REG_DEBUG_BITS]    ip2cpu_debug_reg;
   wire     [`REG_DEBUG_BITS]    cpu2ip_debug_reg; 
   wire     [`REG_RATEBASE_BITS] ratebase_reg;
   wire     [`REG_RATEVALID_BITS] ratevalid_reg;
   wire     [`REG_RATECONFIG_BITS]    rateconfig_reg;


   reg      [`REG_RATEBASE_BITS] time_counter;
   reg      time_expired;
   wire     is_pkt_boundary;
   wire     is_valid_pkt;

   wire clear_counters;
   wire reset_registers;
   wire in_fifo_nearly_full;
   wire in_fifo_empty;
   wire in_fifo_rd_en;
   wire [12:0] data_count;
 
   reg new_packet;


   assign is_pkt_boundary = rateconfig_reg[0];
   assign is_valid_pkt    = rateconfig_reg[4];

uram_fifo #(
	.WIDTH (512+64+128+1),  // 1 to 4096
	.DEPTH (4096)   // 16 to 4194304
) rate_limiter_fifo (
	.clk         (axis_aclk),
	.rst         (~axis_resetn),
	.wr_en       (s_axis_tvalid & ~in_fifo_nearly_full),
	.din         ({s_axis_tlast, s_axis_tuser, s_axis_tkeep, s_axis_tdata}),
	.rd_en       (in_fifo_rd_en),
	.dout        ({m_axis_tlast, m_axis_tuser, m_axis_tkeep, m_axis_tdata}),
	.empty       (in_fifo_empty),
	.full        (),
	.almost_empty(),	 
	.almost_full (in_fifo_nearly_full)
);
//   rate_limiter_fifo
//     //   #( .WIDTH(C_M_AXIS_DATA_WIDTH+C_M_AXIS_TUSER_WIDTH+C_M_AXIS_DATA_WIDTH/8+32+1),
//     //      .MAX_DEPTH_BITS(2))
//      rate_limiter_fifo
//        (// Outputs
//         .dout                           ({m_axis_tlast, m_axis_tuser, m_axis_tkeep, m_axis_tdata}),
//         .full                           (),
//         .almost_full                    (in_fifo_nearly_full),
//         .empty                          (in_fifo_empty),
//         // Inputs
//         .din                            ({s_axis_tlast, s_axis_tuser, s_axis_tkeep, s_axis_tdata}),
//         .wr_en                          (s_axis_tvalid & ~in_fifo_nearly_full),
//         .rd_en                          (in_fifo_rd_en),
//	 .data_count			(data_count),
//         .srst                           (~axis_resetn),
//         .clk                           (axis_aclk));



   assign s_axis_tready = !in_fifo_nearly_full;

 

   // Handle output
   assign in_fifo_rd_en = m_axis_tready && !in_fifo_empty && time_expired;
   assign m_axis_tvalid = !in_fifo_empty && time_expired;


//Registers section
 rate_limiter_cpu_regs 
 #(
   .C_BASE_ADDRESS        (C_BASEADDR),
   .C_S_AXI_DATA_WIDTH (C_S_AXI_DATA_WIDTH),
   .C_S_AXI_ADDR_WIDTH (C_S_AXI_ADDR_WIDTH)
 ) opl_cpu_regs_inst
 (   
   // General ports
    .clk                    (axis_aclk),
    .resetn                 (axis_resetn),
   // AXI Lite ports
    .S_AXI_ACLK             (S_AXI_ACLK),
    .S_AXI_ARESETN          (S_AXI_ARESETN),
    .S_AXI_AWADDR           (S_AXI_AWADDR),
    .S_AXI_AWVALID          (S_AXI_AWVALID),
    .S_AXI_WDATA            (S_AXI_WDATA),
    .S_AXI_WSTRB            (S_AXI_WSTRB),
    .S_AXI_WVALID           (S_AXI_WVALID),
    .S_AXI_BREADY           (S_AXI_BREADY),
    .S_AXI_ARADDR           (S_AXI_ARADDR),
    .S_AXI_ARVALID          (S_AXI_ARVALID),
    .S_AXI_RREADY           (S_AXI_RREADY),
    .S_AXI_ARREADY          (S_AXI_ARREADY),
    .S_AXI_RDATA            (S_AXI_RDATA),
    .S_AXI_RRESP            (S_AXI_RRESP),
    .S_AXI_RVALID           (S_AXI_RVALID),
    .S_AXI_WREADY           (S_AXI_WREADY),
    .S_AXI_BRESP            (S_AXI_BRESP),
    .S_AXI_BVALID           (S_AXI_BVALID),
    .S_AXI_AWREADY          (S_AXI_AWREADY),

   
   // Register ports
   .id_reg          (id_reg),
   .version_reg          (version_reg),
   .reset_reg          (reset_reg),
   .ip2cpu_flip_reg          (ip2cpu_flip_reg),
   .cpu2ip_flip_reg          (cpu2ip_flip_reg),
   .pktin_reg          (pktin_reg),
   .pktin_reg_clear    (pktin_reg_clear),
   .pktout_reg          (pktout_reg),
   .pktout_reg_clear    (pktout_reg_clear),
   .ip2cpu_debug_reg          (ip2cpu_debug_reg),
   .cpu2ip_debug_reg          (cpu2ip_debug_reg),
   .ratebase_reg              (ratebase_reg),
   .ratevalid_reg              (ratevalid_reg),
   .rateconfig_reg             (rateconfig_reg),
   // Global Registers - user can select if to use
   .cpu_resetn_soft(),//software reset, after cpu module
   .resetn_soft    (),//software reset to cpu module (from central reset management)
   .resetn_sync    (resetn_sync)//synchronized reset, use for better timing
);

   assign clear_counters = reset_reg[0];
   assign reset_registers = reset_reg[4];

//a counter used to measure time
always @(posedge axis_aclk)
	if (~resetn_sync | clear_counters) begin
		time_counter <= #1 0;
	end
	else begin
		if (is_pkt_boundary)
			if (is_valid_pkt)
				time_counter <= #1 (ratebase_reg == 0) || (ratevalid_reg == 0) ? 0:
					           !in_fifo_empty & m_axis_tlast & in_fifo_rd_en ? ((time_counter+1 == ratebase_reg) ? 0  : time_counter+1) :
						   time_counter;
			else
				time_counter <= #1 (ratebase_reg == 0) || (ratevalid_reg == 0) ? 0 :
						   (time_counter+1 < ratebase_reg) ? time_counter+1 :
						    (!in_fifo_empty & m_axis_tlast & in_fifo_rd_en) ? time_counter+1 : time_counter ;

		else
			time_counter <= #1 (ratebase_reg == 0) || (ratevalid_reg == 0) || (time_counter+1 == ratebase_reg) ? 0 : 
				            time_counter +1 ; 	
	end

//new packet indicator
always @(posedge axis_aclk)
	if (~resetn_sync) begin
		new_packet <= #1 1'b1;
	end
	else begin
		new_packet <= #1 !in_fifo_empty & m_axis_tlast & in_fifo_rd_en ? 1'b1: in_fifo_empty ? new_packet : 1'b0;
        end	


////registers logic, current logic is just a placeholder for initial compil, required to be changed by the user
always @(posedge axis_aclk)
	if (~resetn_sync | reset_registers) begin
		id_reg <= #1    `REG_ID_DEFAULT;
		version_reg <= #1    `REG_VERSION_DEFAULT;
		ip2cpu_flip_reg <= #1    `REG_FLIP_DEFAULT;
		pktin_reg <= #1    `REG_PKTIN_DEFAULT;
		pktout_reg <= #1    `REG_PKTOUT_DEFAULT;
		ip2cpu_debug_reg <= #1    `REG_DEBUG_DEFAULT;
	end
	else begin
		id_reg <= #1    `REG_ID_DEFAULT;
		version_reg <= #1    `REG_VERSION_DEFAULT;
		ip2cpu_flip_reg <= #1    ~cpu2ip_flip_reg;
		pktin_reg[`REG_PKTIN_WIDTH -2: 0] <= #1  clear_counters | pktin_reg_clear ? 'h0  : pktin_reg[`REG_PKTIN_WIDTH-2:0] + (s_axis_tlast && s_axis_tvalid && s_axis_tready) ;
                pktin_reg[`REG_PKTIN_WIDTH-1] <= #1 clear_counters | pktin_reg_clear ? 1'h0 : pktin_reg_clear ? 'h0  : pktin_reg[`REG_PKTIN_WIDTH-2:0] + (s_axis_tlast && s_axis_tvalid && s_axis_tready) 
                                                     > {(`REG_PKTIN_WIDTH-1){1'b1}} ? 1'b1 : pktin_reg[`REG_PKTIN_WIDTH-1];
                                                               
		pktout_reg [`REG_PKTOUT_WIDTH-2:0]<= #1  clear_counters | pktout_reg_clear ? 'h0  : pktout_reg [`REG_PKTOUT_WIDTH-2:0] + (m_axis_tlast && m_axis_tvalid && m_axis_tready) ;
                pktout_reg [`REG_PKTOUT_WIDTH-1]<= #1  clear_counters | pktout_reg_clear ? 'h0  : pktout_reg [`REG_PKTOUT_WIDTH-2:0] + (m_axis_tlast && m_axis_tvalid && m_axis_tready)  > {(`REG_PKTOUT_WIDTH-1){1'b1}} ?
                                                                1'b1 : pktout_reg [`REG_PKTOUT_WIDTH-1];
		ip2cpu_debug_reg [12:0] <= #1   data_count; //indicate buffer status
                ip2cpu_debug_reg [31:13] <= #1  18'h0;
        end

//Expired time logic
always @(posedge axis_aclk)
	if (~resetn_sync | reset_registers) begin
	   time_expired <= #1 1'b1;
	end
	else begin
	   time_expired <= #1 (ratebase_reg == 0) || (ratevalid_reg == 0) || (ratebase_reg < ratevalid_reg) ? 1'b1 : 
                              time_counter < ratevalid_reg ? 1'b1 : 
			      is_pkt_boundary & !(in_fifo_rd_en & m_axis_tlast) ? 1'b1: 1'b0;
	end
 
endmodule // rate_limiter
